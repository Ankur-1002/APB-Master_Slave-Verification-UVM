package apb_pkg;
    
    //==========================================================================
    // Global Parameters
    //==========================================================================
    `define ADDR_WIDTH = 32;
    `define DATA_WIDTH = 32;  
    `define MEM_DEPTH  = 256;

endpackage: apb_pkg

package master_Pkg;
	`include "uvm_pkg.sv"
	import uvm_pkg::*;
	`include "apb_slave.sv"
	`include "master_tx.sv"
	`include "master_intf.sv"
	`include "master_seq_lib.sv"
	`include "master_mon.sv"
	`include "master_drv.sv"
	`include "master_sqr.sv"
	`include "master_agnt.sv"
	`include "master_env.sv"
	`include "master_test_lib.sv"
endclass

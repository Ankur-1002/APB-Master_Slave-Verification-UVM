class apb_slave_txn extends uvm_sequence_item;

  rand bit 

`include "APB_Define.sv"
`include "apb_intf.sv"
package apb_master_pkg;
 `include "uvm_macros.svh"
  import uvm_pkg::*;
 `include "APB_transaction.sv"
 `include "APB_sequence.sv"
 `include "APB_sequencer.sv"
 `include "APB_driver.sv"
 `include "APB_monitor.sv"
 `include "APB_master_agent.sv"
 `include "apb_env.sv"
 `include "test.sv"

endpackage
